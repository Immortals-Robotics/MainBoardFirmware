module top ( motorin , motorout );
    input[23:0] motorin;
    output[7:0] motorout;
    reg[7:0] motorout;
    always @( motorin )
    begin
        if ( motorin > 3265095 )    motorout <= 0;
        else if ( motorin > 1632547 )   motorout <= 1;
        else if ( motorin > 1088365 )   motorout <= 2;
        else if ( motorin > 816273 )    motorout <= 3;
        else if ( motorin > 653019 )    motorout <= 4;
        else if ( motorin > 544182 )    motorout <= 5;
        else if ( motorin > 466442 )    motorout <= 6;
        else if ( motorin > 408136 )    motorout <= 7;
        else if ( motorin > 362788 )    motorout <= 8;
        else if ( motorin > 326509 )    motorout <= 9;
        else if ( motorin > 296826 )    motorout <= 10;
        else if ( motorin > 272091 )    motorout <= 11;
        else if ( motorin > 251161 )    motorout <= 12;
        else if ( motorin > 233221 )    motorout <= 13;
        else if ( motorin > 217673 )    motorout <= 14;
        else if ( motorin > 204068 )    motorout <= 15;
        else if ( motorin > 192064 )    motorout <= 16;
        else if ( motorin > 181394 )    motorout <= 17;
        else if ( motorin > 171847 )    motorout <= 18;
        else if ( motorin > 163254 )    motorout <= 19;
        else if ( motorin > 155480 )    motorout <= 20;
        else if ( motorin > 148413 )    motorout <= 21;
        else if ( motorin > 141960 )    motorout <= 22;
        else if ( motorin > 136045 )    motorout <= 23;
        else if ( motorin > 130603 )    motorout <= 24;
        else if ( motorin > 125580 )    motorout <= 25;
        else if ( motorin > 120929 )    motorout <= 26;
        else if ( motorin > 116610 )    motorout <= 27;
        else if ( motorin > 112589 )    motorout <= 28;
        else if ( motorin > 108836 )    motorout <= 29;
        else if ( motorin > 105325 )    motorout <= 30;
        else if ( motorin > 102034 )    motorout <= 31;
        else if ( motorin > 98942 ) motorout <= 32;
        else if ( motorin > 96032 ) motorout <= 33;
        else if ( motorin > 93288 ) motorout <= 34;
        else if ( motorin > 90697 ) motorout <= 35;
        else if ( motorin > 88245 ) motorout <= 36;
        else if ( motorin > 85923 ) motorout <= 37;
        else if ( motorin > 83720 ) motorout <= 38;
        else if ( motorin > 81627 ) motorout <= 39;
        else if ( motorin > 79636 ) motorout <= 40;
        else if ( motorin > 77740 ) motorout <= 41;
        else if ( motorin > 75932 ) motorout <= 42;
        else if ( motorin > 74206 ) motorout <= 43;
        else if ( motorin > 72557 ) motorout <= 44;
        else if ( motorin > 70980 ) motorout <= 45;
        else if ( motorin > 69470 ) motorout <= 46;
        else if ( motorin > 68022 ) motorout <= 47;
        else if ( motorin > 66634 ) motorout <= 48;
        else if ( motorin > 65301 ) motorout <= 49;
        else if ( motorin > 64021 ) motorout <= 50;
        else if ( motorin > 62790 ) motorout <= 51;
        else if ( motorin > 61605 ) motorout <= 52;
        else if ( motorin > 60464 ) motorout <= 53;
        else if ( motorin > 59365 ) motorout <= 54;
        else if ( motorin > 58305 ) motorout <= 55;
        else if ( motorin > 57282 ) motorout <= 56;
        else if ( motorin > 56294 ) motorout <= 57;
        else if ( motorin > 55340 ) motorout <= 58;
        else if ( motorin > 54418 ) motorout <= 59;
        else if ( motorin > 53526 ) motorout <= 60;
        else if ( motorin > 52662 ) motorout <= 61;
        else if ( motorin > 51826 ) motorout <= 62;
        else if ( motorin > 51017 ) motorout <= 63;
        else if ( motorin > 50232 ) motorout <= 64;
        else if ( motorin > 49471 ) motorout <= 65;
        else if ( motorin > 48732 ) motorout <= 66;
        else if ( motorin > 48016 ) motorout <= 67;
        else if ( motorin > 47320 ) motorout <= 68;
        else if ( motorin > 46644 ) motorout <= 69;
        else if ( motorin > 45987 ) motorout <= 70;
        else if ( motorin > 45348 ) motorout <= 71;
        else if ( motorin > 44727 ) motorout <= 72;
        else if ( motorin > 44122 ) motorout <= 73;
        else if ( motorin > 43534 ) motorout <= 74;
        else if ( motorin > 42961 ) motorout <= 75;
        else if ( motorin > 42403 ) motorout <= 76;
        else if ( motorin > 41860 ) motorout <= 77;
        else if ( motorin > 41330 ) motorout <= 78;
        else if ( motorin > 40813 ) motorout <= 79;
        else if ( motorin > 40309 ) motorout <= 80;
        else if ( motorin > 39818 ) motorout <= 81;
        else if ( motorin > 39338 ) motorout <= 82;
        else if ( motorin > 38870 ) motorout <= 83;
        else if ( motorin > 38412 ) motorout <= 84;
        else if ( motorin > 37966 ) motorout <= 85;
        else if ( motorin > 37529 ) motorout <= 86;
        else if ( motorin > 37103 ) motorout <= 87;
        else if ( motorin > 36686 ) motorout <= 88;
        else if ( motorin > 36278 ) motorout <= 89;
        else if ( motorin > 35880 ) motorout <= 90;
        else if ( motorin > 35490 ) motorout <= 91;
        else if ( motorin > 35108 ) motorout <= 92;
        else if ( motorin > 34735 ) motorout <= 93;
        else if ( motorin > 34369 ) motorout <= 94;
        else if ( motorin > 34011 ) motorout <= 95;
        else if ( motorin > 33660 ) motorout <= 96;
        else if ( motorin > 33317 ) motorout <= 97;
        else if ( motorin > 32980 ) motorout <= 98;
        else if ( motorin > 32650 ) motorout <= 99;
        else if ( motorin > 32327 ) motorout <= 100;
        else if ( motorin > 32010 ) motorout <= 101;
        else if ( motorin > 31699 ) motorout <= 102;
        else if ( motorin > 31395 ) motorout <= 103;
        else if ( motorin > 31096 ) motorout <= 104;
        else if ( motorin > 30802 ) motorout <= 105;
        else if ( motorin > 30514 ) motorout <= 106;
        else if ( motorin > 30232 ) motorout <= 107;
        else if ( motorin > 29955 ) motorout <= 108;
        else if ( motorin > 29682 ) motorout <= 109;
        else if ( motorin > 29415 ) motorout <= 110;
        else if ( motorin > 29152 ) motorout <= 111;
        else if ( motorin > 28894 ) motorout <= 112;
        else if ( motorin > 28641 ) motorout <= 113;
        else if ( motorin > 28392 ) motorout <= 114;
        else if ( motorin > 28147 ) motorout <= 115;
        else if ( motorin > 27906 ) motorout <= 116;
        else if ( motorin > 27670 ) motorout <= 117;
        else if ( motorin > 27437 ) motorout <= 118;
        else if ( motorin > 27209 ) motorout <= 119;
        else if ( motorin > 26984 ) motorout <= 120;
        else if ( motorin > 26763 ) motorout <= 121;
        else if ( motorin > 26545 ) motorout <= 122;
        else if ( motorin > 26331 ) motorout <= 123;
        else if ( motorin > 26120 ) motorout <= 124;
        else if ( motorin > 25913 ) motorout <= 125;
        else if ( motorin > 25709 ) motorout <= 126;
        else if ( motorin > 25508 ) motorout <= 127;
        else if ( motorin > 25310 ) motorout <= 128;
        else if ( motorin > 25116 ) motorout <= 129;
        else if ( motorin > 24924 ) motorout <= 130;
        else if ( motorin > 24735 ) motorout <= 131;
        else if ( motorin > 24549 ) motorout <= 132;
        else if ( motorin > 24366 ) motorout <= 133;
        else if ( motorin > 24185 ) motorout <= 134;
        else if ( motorin > 24008 ) motorout <= 135;
        else if ( motorin > 23832 ) motorout <= 136;
        else if ( motorin > 23660 ) motorout <= 137;
        else if ( motorin > 23489 ) motorout <= 138;
        else if ( motorin > 23322 ) motorout <= 139;
        else if ( motorin > 23156 ) motorout <= 140;
        else if ( motorin > 22993 ) motorout <= 141;
        else if ( motorin > 22832 ) motorout <= 142;
        else if ( motorin > 22674 ) motorout <= 143;
        else if ( motorin > 22517 ) motorout <= 144;
        else if ( motorin > 22363 ) motorout <= 145;
        else if ( motorin > 22211 ) motorout <= 146;
        else if ( motorin > 22061 ) motorout <= 147;
        else if ( motorin > 21913 ) motorout <= 148;
        else if ( motorin > 21767 ) motorout <= 149;
        else if ( motorin > 21623 ) motorout <= 150;
        else if ( motorin > 21480 ) motorout <= 151;
        else if ( motorin > 21340 ) motorout <= 152;
        else if ( motorin > 21201 ) motorout <= 153;
        else if ( motorin > 21065 ) motorout <= 154;
        else if ( motorin > 20930 ) motorout <= 155;
        else if ( motorin > 20796 ) motorout <= 156;
        else if ( motorin > 20665 ) motorout <= 157;
        else if ( motorin > 20535 ) motorout <= 158;
        else if ( motorin > 20406 ) motorout <= 159;
        else if ( motorin > 20280 ) motorout <= 160;
        else if ( motorin > 20154 ) motorout <= 161;
        else if ( motorin > 20031 ) motorout <= 162;
        else if ( motorin > 19909 ) motorout <= 163;
        else if ( motorin > 19788 ) motorout <= 164;
        else if ( motorin > 19669 ) motorout <= 165;
        else if ( motorin > 19551 ) motorout <= 166;
        else if ( motorin > 19435 ) motorout <= 167;
        else if ( motorin > 19320 ) motorout <= 168;
        else if ( motorin > 19206 ) motorout <= 169;
        else if ( motorin > 19094 ) motorout <= 170;
        else if ( motorin > 18983 ) motorout <= 171;
        else if ( motorin > 18873 ) motorout <= 172;
        else if ( motorin > 18764 ) motorout <= 173;
        else if ( motorin > 18657 ) motorout <= 174;
        else if ( motorin > 18551 ) motorout <= 175;
        else if ( motorin > 18446 ) motorout <= 176;
        else if ( motorin > 18343 ) motorout <= 177;
        else if ( motorin > 18240 ) motorout <= 178;
        else if ( motorin > 18139 ) motorout <= 179;
        else if ( motorin > 18039 ) motorout <= 180;
        else if ( motorin > 17940 ) motorout <= 181;
        else if ( motorin > 17842 ) motorout <= 182;
        else if ( motorin > 17745 ) motorout <= 183;
        else if ( motorin > 17649 ) motorout <= 184;
        else if ( motorin > 17554 ) motorout <= 185;
        else if ( motorin > 17460 ) motorout <= 186;
        else if ( motorin > 17367 ) motorout <= 187;
        else if ( motorin > 17275 ) motorout <= 188;
        else if ( motorin > 17184 ) motorout <= 189;
        else if ( motorin > 17094 ) motorout <= 190;
        else if ( motorin > 17005 ) motorout <= 191;
        else if ( motorin > 16917 ) motorout <= 192;
        else if ( motorin > 16830 ) motorout <= 193;
        else if ( motorin > 16744 ) motorout <= 194;
        else if ( motorin > 16658 ) motorout <= 195;
        else if ( motorin > 16574 ) motorout <= 196;
        else if ( motorin > 16490 ) motorout <= 197;
        else if ( motorin > 16407 ) motorout <= 198;
        else if ( motorin > 16325 ) motorout <= 199;
        else if ( motorin > 16244 ) motorout <= 200;
        else if ( motorin > 16163 ) motorout <= 201;
        else if ( motorin > 16084 ) motorout <= 202;
        else if ( motorin > 16005 ) motorout <= 203;
        else if ( motorin > 15927 ) motorout <= 204;
        else if ( motorin > 15849 ) motorout <= 205;
        else if ( motorin > 15773 ) motorout <= 206;
        else if ( motorin > 15697 ) motorout <= 207;
        else if ( motorin > 15622 ) motorout <= 208;
        else if ( motorin > 15548 ) motorout <= 209;
        else if ( motorin > 15474 ) motorout <= 210;
        else if ( motorin > 15401 ) motorout <= 211;
        else if ( motorin > 15329 ) motorout <= 212;
        else if ( motorin > 15257 ) motorout <= 213;
        else if ( motorin > 15186 ) motorout <= 214;
        else if ( motorin > 15116 ) motorout <= 215;
        else if ( motorin > 15046 ) motorout <= 216;
        else if ( motorin > 14977 ) motorout <= 217;
        else if ( motorin > 14909 ) motorout <= 218;
        else if ( motorin > 14841 ) motorout <= 219;
        else if ( motorin > 14774 ) motorout <= 220;
        else if ( motorin > 14707 ) motorout <= 221;
        else if ( motorin > 14641 ) motorout <= 222;
        else if ( motorin > 14576 ) motorout <= 223;
        else if ( motorin > 14511 ) motorout <= 224;
        else if ( motorin > 14447 ) motorout <= 225;
        else if ( motorin > 14383 ) motorout <= 226;
        else if ( motorin > 14320 ) motorout <= 227;
        else if ( motorin > 14258 ) motorout <= 228;
        else if ( motorin > 14196 ) motorout <= 229;
        else if ( motorin > 14134 ) motorout <= 230;
        else if ( motorin > 14073 ) motorout <= 231;
        else if ( motorin > 14013 ) motorout <= 232;
        else if ( motorin > 13953 ) motorout <= 233;
        else if ( motorin > 13894 ) motorout <= 234;
        else if ( motorin > 13835 ) motorout <= 235;
        else if ( motorin > 13776 ) motorout <= 236;
        else if ( motorin > 13718 ) motorout <= 237;
        else if ( motorin > 13661 ) motorout <= 238;
        else if ( motorin > 13604 ) motorout <= 239;
        else if ( motorin > 13548 ) motorout <= 240;
        else if ( motorin > 13492 ) motorout <= 241;
        else if ( motorin > 13436 ) motorout <= 242;
        else if ( motorin > 13381 ) motorout <= 243;
        else if ( motorin > 13326 ) motorout <= 244;
        else if ( motorin > 13272 ) motorout <= 245;
        else if ( motorin > 13219 ) motorout <= 246;
        else if ( motorin > 13165 ) motorout <= 247;
        else if ( motorin > 13112 ) motorout <= 248;
        else if ( motorin > 13060 ) motorout <= 249;
        else if ( motorin > 13008 ) motorout <= 250;
        else if ( motorin > 12956 ) motorout <= 251;
        else if ( motorin > 12905 ) motorout <= 252;
        else if ( motorin > 12854 ) motorout <= 253;
        else if ( motorin > 12804 ) motorout <= 254;
        else    motorout <= 255 ;
    end
endmodule
